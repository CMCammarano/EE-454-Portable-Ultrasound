`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   20:12:24 10/05/2015
// Design Name:   quickhull.v
// 
////////////////////////////////////////////////////////////////////////////////

module m_quickhull_tb;

	// Inputs
	reg CLK100MHZ;
	reg CPU_RESETN;
	reg [4095:0] points;
	reg [7:0] SS;

	// Outputs
	wire [4095:0] convexPoints;
	wire [7:0] convexSetSize;
	wire [7:0] positiveCrossCount;
	wire [15:0] crossValue;
	wire [15:0] lnIndex;
	wire [7:0] ptCount;
	wire [31:0] currLine;
	wire [15:0] currPoint;
	wire [15:0] furthest;

	wire QINITIAL, QFIND_MAX, QFIND_MIN, QHULL_START, QCROSS, QHULL_RECURSE, QEND;
	// File
	integer file_results;

	// Parameters
	parameter CLK_PERIOD = 20;

	// Instantiate the Unit Under Test (UUT)
	m_port_ultra_quickhull_processor UUT(
		//Inputs
		.CLK100MHZ(CLK100MHZ),
		.CPU_RESETN(CPU_RESETN),
		.SS(SS),
		.points(points),
		//Outputs
		.convexPoints(convexPoints),
		.convexSetSizeOutput(convexSetSize),
		.positiveCrossCountOutput(positiveCrossCount),
		.crossValueOutput(crossValue),
		.lnIndexOutput(lnIndex),
		.ptCountOutput(ptCount),
		.currentLineOutput(currLine),
		.currentPointOutput(currPoint),
		.furthestOutput(furthest),
		.QINITIAL(QINITIAL),
		.QFIND_MAX(QFIND_MAX),
		.QFIND_MIN(QFIND_MIN),
		.QHULL_START(QHULL_START),
		.QCROSS(QCROSS),
		.QHULL_RECURSE(QHULL_RECURSE),
		.QEND(QEND)
	);


	initial begin : CLOCK_GENERATOR
		CLK100MHZ = 0;
		
		forever begin
			# (CLK_PERIOD / 2) CLK100MHZ = ~CLK100MHZ;
		end
	end	
		
	integer counter;
	
	initial begin : STIMULUS
		
		//file_results = $fopen("output_results.txt", "w");

		// Initialize Inputs
		// === Small input: 15 points ===
		CLK100MHZ = 0;
		SS = 15;
		CPU_RESETN = 1;
		points = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000101000010000000001100000111000001110000100100000111000001000000001000000101000001010000000100000100000001100000010100000011000001000000001000000100000001010000010100000110000000110000010000001100000010010000101100000001;
		
		for (counter = 0; counter < convexSetSize; counter = counter + 1) begin
			//$fwrite(file_results, " %h", convexPoints[(16*counter)-1 +: (16*counter)]);
			//$write(file_results, " %h", convexPoints[(16*counter)-1 +: (16*counter)]);
		end


		// Wait for global reset to finish
		#100;
				
		// Generate a reset
		CPU_RESETN = 0;	#20;
		CPU_RESETN = 1;	#20;
		
		// Give a long time for machine to finish
		#500000;
		
		/*
		//$fwrite(file_results, "Points:     ");
		$write("Points:     ");
		
		// Wait for global reset to finish
		#100;

		// === Medium input: 50 points ===
		//Input next test
		SS = 50;
		points = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010011011010100101110011101110110011011001000001010100010010010001101100111110010111010110011010000000100001011110000001011110010001001110010010010110101110010111100001101101101000110010011101110001100000011111000011111010110100111010100000110110110110111010110010111011010011101010100001110101101101001110101101010101011111100100011100010100101111110011111101000110100001010011010101110001110011101110110100001000010101111000101001000101100011100000000010101011001010110101101011000100010010111001101011011110110010010010101000101110001100000000101100001110010010111001000011111010001001100100000100010001110101010010110111010001011111011110111111000111110011011001001001010001010000010101001100011100000101000001100011011011000111000101110001110011101001010110101011001011011011010100100011110000011;

		for (counter = 0; counter < convexSetSize; counter = counter + 1) begin
			//$fwrite(file_results, " %h", convexPoints[(16*counter)-1 +: (16*counter)]);
			//$write(file_results, " %h", convexPoints[(16*counter)-1 +: (16*counter)]);
		end


		// Wait for global reset to finish
		#100;
				
		// Generate a reset
		CPU_RESETN = 0;	#20;
		CPU_RESETN = 1;	#20;
		
		// Give a long time for machine to finish
		#5000;
		
		//$fwrite(file_results, "Points:     ");
		$write("Points:     ");
		
		// Wait for global reset to finish
		#100;

		// === Max input: 256 points ===
		// Input next test
		SS = 255;
		points =  4096'b0101110111110101111110100000100001100000111110100110001101001011011010000010110001110001100000011000011111001101011101100001010100010100000010111000111100011000101110101110011101000100101010110010100100010111100111000110011000010010000110010111111010000011000100000001110111101100001110001100001110000100010110111110100110011011011000000100010110001001001011100001111110100101101001101101000010010001011110001010100000100001010111011101110011000011001000001100011001111010111000110010000101111101110110110101000000011011001100100111110010101101100011111010010101001001010010110111011111100100100100001111110011111001100010000110100101100011101010001010001011000110010000010110101110001011011001001000100011100011000100110011000101111010010100010100101110100010011000111011011001011011011100000011010001100101110111101111111100101010101101001100011010111000100010101110101010111100111100000010011101101011101110000100011011011010110111000101100111100001111110101110000111010110111111011101010100100010011001010001111000110110010011110110010110000100001000010001110100110110111101000000000001011010110000111101100001111010000001100111111010101110111010110010110010110100110100010101000001010000011110001100101001010001011011100100110111001011010000100011001000001001000011101010010010100011010100001110100011100000000101101111000110000110000001000100100110000010010001100101000011001111011010110010111010100110111101000101000111101111001010010011101100110111010010111110001111011010000000010011111110100010100010010011010111010101101110000100000010110000111000110111000011111000001011001101100010110110100101010100111010110100000011010000100100110100101001100100010110101000010010110011111100011011110001001101001110001110000110011000001101001010011011011110000000100001001010100010001101100101111011110011001111001111001011110011110101001001011011011011111011110000100110011110101101010111010011101110011011101010111101110010111101110101110010011110001000000111010010100001110001001001010001010100110001110110001011010001110111110011000100111000110111001111100100111110000100000111000101110110111011110101100001000001011111000100001100000111010110000010010011011101100100111000001011011100011010111111001011010101101000011110000111100001001010010001111110011001111011111011001010111111111110111101101000100111110101011111111001000111110011000111110110000000101011010111101010101101101000111110100000000001101111100110101110011010001000111010010101110101101001010000011110111101000111000011000001110101100010100110001001000000100001010000010101110011011001110110011010100110001001000001001101010101111011110111011011011111111010110100011101011000000011010010001011100000000000100101000011101001010000000001110001101111100001000010100100001010111001010100010101100100101001111010010000000010011111000010101011101001111010011010110110100010101010100111011111001000101000010110100111000010000001010001011001011000100011111001010010000011100010001011001001100000110100001011000110100011001101000110110000001001101000101111111111011010101100101110111010111010001110001101001011110010111001000101100010000011101011110011001001100110011100001010000111100011001110001101101010011110100000100011100001101111101010101111110100101111100001110000101000001001111110010010101000000001010001001011111000011001110110010101001011000101101011100101110110111001110010110011000101000011001000110010001011110101000100110001110110011111001000111010111110001000010101111111010011111011111111010110001010000100011001101000011000111000110010010001100101011100001100100010011111100000111101110011101101100000000110110100001010111111010001011110011000101001011100001100001111001010010010001011000001000100101010011100010001101010001110001110000001010000100111011100111100100110101101001101111111010001110100100100001101101010111110000010011010010101010100010101011010111101010001100011001001111011010111110011110011110001110100110100001010111011000111011001101110100101111100001100100011001010111101111000001001000010110101010101110011000011101110001000110011100110001110101011110000001001100101100101010101011111110101011010;

		for (counter = 0; counter < convexSetSize; counter = counter + 1) begin
			//$fwrite(file_results, " %h", convexPoints[(16*counter)-1 +: (16*counter)]);
			//$write(file_results, " %h", convexPoints[(16*counter)-1 +: (16*counter)]);
		end


		// Wait for global reset to finish
		#100;
				
		// Generate a reset
		CPU_RESETN = 0;	#20;
		CPU_RESETN = 1;	#20;
		
		// Give a long time for machine to finish
		#10000;
		
		//$fwrite(file_results, "Points:     ");
		$write("Points:     ");
		*/
		// Wait for global reset to finish
		#100;

	$fclose (file_results);	 

	end
		  
endmodule

