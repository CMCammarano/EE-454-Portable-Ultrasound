`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   20:12:24 10/05/2015
// Design Name:   quickhull.v
// 
////////////////////////////////////////////////////////////////////////////////

module m_port_ultra_tb;

	// Inputs
	reg CLK100MHZ;
	reg CPU_RESETN;
	reg BTNC;
	reg [32767:0] convexCloud;

	// Outputs
	wire [4095:0] convexHull1;
	wire [4095:0] convexHull2;
	wire [4095:0] convexHull3;
	wire [4095:0] convexHull4;
	wire [4095:0] convexHull5;
	wire [4095:0] convexHull6;
	wire [4095:0] convexHull7;
	wire [4095:0] convexHull8;
	wire [8:0] convexHullSize1;
	wire [8:0] convexHullSize2;
	wire [8:0] convexHullSize3;
	wire [8:0] convexHullSize4;
	wire [8:0] convexHullSize5;
	wire [8:0] convexHullSize6;
	wire [8:0] convexHullSize7;
	wire [8:0] convexHullSize8;
	wire processorDone1;
	wire processorDone2;
	wire processorDone3;
	wire processorDone4;
	wire processorDone5;
	wire processorDone6;
	wire processorDone7;
	wire processorDone8;
	wire QINIT, QPULSE, QDIVIDE, QCONVEX_HULL, QDISPLAY;

	// Parameters
	parameter CLK_PERIOD = 20;

	// Instantiate the Unit Under Test (UUT)
	m_port_ultra UUT(
		.clk (CLK100MHZ),
		.reset_n (CPU_RESETN),
		.ack (BTNC),
		.convexCloud (convexCloud),
		.convexHull1 (convexHull1),
		.convexHull2 (convexHull2),
		.convexHull3 (convexHull3),
		.convexHull4 (convexHull4),
		.convexHull5 (convexHull5),
		.convexHull6 (convexHull6),
		.convexHull7 (convexHull7),
		.convexHull8 (convexHull8),
		.convexHullSize1 (convexHullSize1),
		.convexHullSize2 (convexHullSize2),
		.convexHullSize3 (convexHullSize3),
		.convexHullSize4 (convexHullSize4),
		.convexHullSize5 (convexHullSize5),
		.convexHullSize6 (convexHullSize6),
		.convexHullSize7 (convexHullSize7),
		.convexHullSize8 (convexHullSize8),
		.processorDone1 (processorDone1),
		.processorDone2 (processorDone2),
		.processorDone3 (processorDone3),
		.processorDone4 (processorDone4),
		.processorDone5 (processorDone5),
		.processorDone6 (processorDone6),
		.processorDone7 (processorDone7),
		.processorDone8 (processorDone8),
		.QINIT (QINIT),
		.QPULSE (QPULSE),
		.QDIVIDE (QDIVIDE),
		.QCONVEX_HULL (QCONVEX_HULL),
		.QDISPLAY (QDISPLAY)
	);


	initial begin : CLOCK_GENERATOR
		CLK100MHZ = 0;
		
		forever begin
			# (CLK_PERIOD / 2) CLK100MHZ = ~CLK100MHZ;
		end
	end	
		
	integer counter;
	
	initial begin : STIMULUS
		
		// 256 per processor, 64
		convexCloud = 32768'b00001111000000000010110000101001001010100011000000000110000001110010110000011010001111100000110000100011000111000010001000001000000011000011110000110101001110000011111000110100001101110011011100011011001111100000110100111001000001010010100100101010000101010001011100001000001110100000001100101111000101100010011000011011001100010011101000011001000011100010001000111000000000100011011000101111000001100001010100010001001011110011011100011001001010000011101000101111001101010011110000011101000101100010111000101110000000110011011100111001001011100000111000010000000111000011111000101001001101000000110100001110001110110001110100111000001000000010100100010000000111110010010100000111001010100010000100101001000001100001000000101111000000100010011100101010001100010010010100010111001001100001001000111000000011000011110000000001001100010001001100100111000111110010001100111000000001110011000000010001000001000010010000000100001000100001011100011100000001110001001100001100001000100001100000110101001000100011010000111000001101110011110000101111001010110011011000101101000010000010001100101101000101000011000000100000000100110010100000110000001101010001001000011001001000010010100100010010001101100001001000011010000011110011011000111000000110010001101000001010001000100000010100100010000101000001000000000101001110110000111100100110000001110010001100001110001011110010100000010010001100100011101100011110001110000010001000111100000001100001100000000011001011000000101100110011001100000001111100101110000011110001011100110011000000000001111000101110000000010011011100101001001100000001001000010101001101000000010100110101001110000011110000111010001010010001010100011100000010100010101000111001000100110010100000110100000010110001101100111011000101000001011000000010000010000011011000010110001001000000101000110001000010110001000000111100001101000001100100111101001000100000100000001110001010100011101000100110000101010000001100011100001110110011111100100101000101000010011100000100001001110010011000110001000110110001100000000001000010110011111100101011000010010000000100110000000110100011101000000100001000110000111000111100001010000000011000110000001000000001001000110101000011000000110100111010000001110000000100010000001001110001111100111010001101100001011000010110000010010010000100000011001111110010111100100111000000010011000000001011001101110010001100001001001011000000111000110111000110100011110100110111000001010011011000010011001001100000110000101000001011010000111000101000000110010001100100101011001011010010111000101111000101000000100100100101000011000010010000110000001001010001101100001100000001000011010100000100000000000001100100101111000000000010001100100100000100010000101000001111001110100001011000001111000111110000111000100001001011110011101100110001001110010010001000000011000100000001110100100111000010010010100100110001000111000000011000110000001010100010010100101110001111110011110100000101000001010011101100001011001101010011001100011001000000100001110000000010001010000011011000100110000001000000100000010011001010010010011000010011001011010010010100110110000110100001101100110011000011010000011000010111000100010000001100000110000110110000110000101110001101110010100000111011000101100001110100000101000010100011001000000010000011000010001000011000000110010000100000111110000101100000101100111100001100110000011000000101001110110001111100110010001001110010000100010101001011000010010000110100001010010011110000010001000100000010001100111110001000000010010000111100001100000010011100101010000010110001011100010011000110010001100000110000000000100011001000011101001011000000010000001001001110000001110000110011001110110011100100101001001010000011100100010001001110000000010100001011000010010010110000010101001010100001001000011110001111010011010100010000001001100001001100011000001000100001010000011011000000010001111100100110000010000011001100010111001100100010101000001010001111000010011000110001001010010001110000001000001101110011000100000000001001000000111100110000000100110010111100011111000101000011101100110111001111100010110000000111001111000000101000110011001110010011000100101001000101100000001100100101000011000010101100000011000010110011110000010011001110000010110100000100000010000010011000000101000100100011011100100000000001110000010000111110000001110001100100000101000111010010110100011010001010010000011000111010001100000010111000001001001010010001000000111001000011110010110100001011000010110010101100100011000100010010010000110101000111010000110000111000001100110010011100011101000000000011110000011100000000000011000100010000001011100001001000111101001111000001110100000100000000010001101100100001001100010010011000010000000011010000011000011110001100110000110100000011000111010010000000000101000110100010001100010000000011010011010000011000001010000010110100010011000101110001101100001101001111110011101000011010001000000000101100011000001010000010100100001101000110010000100100101111001111010000011100010000000001010011010000001100001111000010110000000110000100000010011000100011001110000010101000010011000000010000010000101010000001100001110000010010001100010011011000100111000100100010001000111101001001010010101100111001001001110011000000010100000110110011011100000001001001110000001000011011001010010011000100010011000001000010000100001110000010100001011000101101000011100000101000011110000100110001010000000010001011100001000000100011000010000011011100110101000000000000110100000011001101100011001000010011000111110000010000110101000101010010010000010010000100010000111100111011001011000011111000010000000100100000110100110010001011110000110100110001000000110001000000111101001001100011001000110111000011000011100000101000001110100000011100000000000001010010110100111111001111110011010000100110001001010000010100111101000101100011101000011110000000000010111000101001001000010011010000001011001111000010111100001110000011110010111000100001000010010010000000101111001101110010101100000101001111100000111000110011001000010000011000100111001111100000001100110001000110100011001000101010001011100000000000001011000011100010010100101000001101100000011000100001001000000001011100101111000001000000101000000010001000100010110100110100000100000010110000100010001100000011111100110110001101110011001000011010000011100011001000100101001101100011101100111100000001110010110100101001001110110000011100110010000101110000011000000101001000110011001100100110000101010011111000110111000101110000000000101101000101110000101100110010001010010001001000000010000110110001101100110000000001100001111000001001001101110011100100111001001100010000001100001110001101100000110100110001001001100000111000001001000010010001000000000001001000110000001100111011000111100001011000001010000100110001111000100100000011110000100000101100000101110000000100011011000110000010010000011110001100000011011000100100000110110011001100000011001100100001010000100100001110100011010100100000000110010010000000011001000110110001011100111110001110010001010000100011000010000001010000110011000011110001010000101011000010000001100000101100001001000010100100001111001010110011110000011010001101110001011100100100000011000000001100100001001111110010110100100110001101000011110100100011000100100011110100111011001001000001010000001110001010110001110000101001000011110011111100001101001111000011010100011100001110110010101100010010001000000010011000010111000001110001011000001110001100000011010100011100000000010010110100010000001100100000011100001001001000110010001000100100001010110000110100010100001011010001001100001001001101110001101100011001001100010000011100010110001001000011100100011100001110110001100000100000001001110000101100001101000000010000100000010001001001010010001000001001001111110010001000001000001111000010101100110110000100010010001000100010000001110011000000010111001000000000101100101000000011100001111000111001000111010010110000000000000110100010011000111001000001000000101100011100000001100001001100011001000101100011011000111111001001010011011100111011001001000000000000010100001010000000111000100011000111100010100000010000000110110000011000111011001111000000111000111100000000110001100000000011001100010011011100100000001100100010111000100011000001000000011100101000001110110011001000100110000111010000001000011000000110100011110000011000001110100001010100000100000010010000100100001111000000100000110100000000000111110011101100000011001010010010111000000000001001100001001000111101000000010011110000011111000111010010101000011010000110100011011000100000000011010010000100001000000011100001100000100010001001010011010100111011000100110000111100110000000100010011001000011010001000110010100000110001000000010010001100111111000000000000101000000100001111000010110100001011000010110001101100100011001111110010001100101010001011100001011000011010000111110000100000111111000010010011010000111000001001010001011100000010001111100000001100010100001101100000011100001111000110100000001000110111000111000000010000010010000010010011111000111111000101010010111100101010001000100001110100110001001000010011011100000011001010000010011100100111000110100000110100011000001100100010011000101011000001100010010000110000000000010011110100010110000100110001001100100011001111000000010000101000001100000000001000001000000011010001010000001000001011100001111100000100001101110001110000011000001101100000010000000111001110110010011000010111000100000010101000001010001101100010011000010111000110000000011000101100001010100001001000100001001110010000011100010110001001100011101000111100001101100010111000101001000111010000000000010100000111000001000000101000001101000001101100101001000001100001011000100000000111100011010100101100000101010000010000010101000010110010100100111001001000010000001000101010000111000000110100101000000110100001111100001000000001100000100100010011000010000001000100110010001011000001010100000110001100110000001100011111001110000011000100000000001000010001000100111101001010010010001000101010001100110010110100101101001111010011000100101111000010110010000000011011000100010011110100000011001011100010000100010111001101100011000100000100000101010000011000110010001100110001001100111000000101000010000000100001001100100010000100111000000011000001001000101111000001110010101100001101001111110010111000111111000001100010110100100110001101000011111000110010000001010001110100011000001001100000010000100110001100010011011000000010001101010010011000000100000011010001101100111110001111000011110000101101000101110010110000011110001101000000000100001111001101010001111100111101001111000001011100111111000001100010010100001111000001000011101000110101000111000010101000111101000110010010001100000010001011010011101100110010000100010011101000001110000110110001000100001100001110000011111000000111000000010001100100110110000011110010001000111101001110110011111000011001000001010000001100000110000101110000111000111101000010010000011100011101000000000000101000101001000010000001001100111010000111010000000100100000001011000000001100111010001000100001010000010100000011110011001000101111000001010001101100001111001100110010001000000111000111000000010100100110000101000000110000101001000110100000011100101001000111010010011000110010000101010001000100001010000001000011101000001111001100110001111100011000001011110010100100010110001111100011111100011100000101110001111000100000000010110001100100110100000011100000010100111010001110110010011100001011000011110011011100000011000001110010111100011111001010010011110000001000000000110000110100011010001001100000100100111001001101100000101100010011000110010000000000010010001110000010101000110011001010010010010000101000001110010000001000101110001010110000111000111010000110010010110100010101000000100001010000101110001111110001001100110100000110110010000000100001000010010000011100011101001111000000011100010111000000110010110000111101000111010010101000000110001000110011011000110110000000010010001000011110001111110000000000100111000110110001001000111111000001000010011100111011000000010000110100001111001110010001101100111000000010100000000000010110001000100010100100110100000010010000101100101010000100000000100000000010001010110000000000111011001111000011000100101011001000000011010000100100001110000001010100110011000011100001110100101011000000110010100000010001001111010001100100001110000101000000010000111100001101110010000000000100001011000001100100010001000011100011111100001001000010110011010100000100001010110000100100011011000110010010010100010000000100110011101000110011000001000011011100001001000111010001111000111110000111000001100000100110001011100000000100111000001110000000001000010010001110110010100000000001000110110001101100110111001000000000010000111111001101000000110100000101001110010011110000001010001000110010100100110100001001100011001100111001000010110011010000000010001010100001010000100011001111010010111100110000001011110011111100101011000111010010010100111100000010110011110100011000001101100011011100101000001001010010000000111011001111100011010000111101000101000001110100011001000000100001111000010101000100010001010100001011000001010000101000111000000110100010001100011111001111000001011100101100000100100010101000001101000011100000100100100010001111000010000100110011000111000000000100011011000100010001110000100111000101100010110000011011001001000000010000001111000000000001100000100010000010010000100000101100000101010010011000000110001110000001010100100010001010000000110100000001001001000000110100111101001011010010110100110011001100100010111100110110000110100000101100111011001100010010010100010110000111010010111000011100000101000001111100001100001111110000010100111111000110000010000100011011000101110001101100111100001011110011110100010000000001110011100000101110001100110010011000001100000001100011111000110001000110010011100000001100000100100000101100001001001101000000100000000101000100010011100100101110001000000010100100000101000110110001001100000101000011110011111100000001001101010001001000110000001010000000011000000000001011010010110100011111000011100001100000100000000100100001100100111110000100110001001000110110001000110010100000000100001011100000001100101011000000010000101000001110001100000001011100001101000010010000000100000100000110010000110000001111000001110001001100101111001011000010001100101111001101010010010000101000001011000011101100001000000111110001001100011000000111110000101100011100000100100011011100010100001110100000011100010110001101000000010000110000001011100000011100000010000100100001100000000010001100010011100000000101001110000001100000000000000000110011011000000000001110110000101100001100000001110011000100011000000010010010101100011111001111010001000100000110000001010001000100110101001011000010110100101010001100100000011000111111001101000011001000011000001111000010010100010011001101100011010100100011000100110010010100111110001101100010110000101110000110000000011100110000000100010010100000001001000001010000010100111110000010110001111000111101000111000010001000110001000000110010000100101101000000110011000100111101001101100010110000010011001100100011000100010001000000110000011000001110001010010010010100000000000000010000001100111001000100110011001100011111000111010011111000010011000100110010010000011111000011010011100000111101000100010011111100000101001110110000001000100111000011010000011100110010001000000010010100000000000100010010000000010010001101010000110000000011001100100010111100001111000001110001001100010000000110100011100100011011000011110010110000001010000101010001101000111110001010110000100000111001000111010001010000000011000101010001011100011010001110110010000000110100000100100000000100000001001111110001110100100000000001100011100100010100000110110011011000010111000110100001010000011011001001000010111100001001000011010011111100111000001110000010011000100111000000110011000100000110001111100010001100000011001100000011011000001111001100010000001000001111001011010011001100000100000110000000001000101000001011100001011100100101000001110001011000100001001011010001010100100010001101110010101000100101000101110011001000011100000001000001000000011110001101000001100000101101001100010010111000001001000110110000011100100001000001010001111000000111001010100000000000010100001101110001001100000110001101100001001000110111000000000010101100010100000011110000011000000001001111000000011000000111000110100010000000011101000001010011001100010100000000110001100000110011001011100010011100101111000101100000110000000000001100010010011100111110001110010001111100111110001101100011000100000101000010010001001100100110001000000010011100010110001111010010111000010100000011000000111100100100000001100000001000110111001010100011100100101100000100000010000100101100001111110011111100010111000011000001000000111110000110100000001100010010001101100011001100110011001001010010010000000010001110110010000100000111001110110000100000000111001010010000110000110101000001110010001000011100001000110001001000111110001110010001011000010101001000000010111000011011000111010000101000100101000110010011111100111110000110110000001000001110001000010001000000010110001000100000001000000011001010110010100100010110000101110011101100000101000000100000011100011011001111100011110100001000000000100011110000111000000111000010001000010000001111010011100100001110001001110010010000110110001011110001111100101110000001000011000000010111000010010011001000110000001111100001011100110100001110010000111000011000000110100010100000010111000101000011000100000011001000010010000100011101000111010000101000110100000000100001001000010111000101000011101100100010000110100001111000101111001110100010010100000000000111110001001100011101001101110001100000100011001001110001001100011110000111100001110000011011001111110001000100000101000110110000010000100111000100100010100000101111000001010011001000001101000011000001110100111000001011000000001000110000001111100001100000110000001110000001001000010101001010110001001000111100000010110010100100010000000111010000000000001111000110100010111000100000000110000011100100110100000011100001011100100110001110110011100000110110000000000011000100111001001101110011001000011100001011100000100100000011001001100010000100011001001011000010000000110101000111100001101000011101001000010001001100111011000001010000111000110000001101100001011000101100001101110011100000110111001111000010101000010110000000100001001000110001000101100001001100011100000001000010001000010000000100010011101100010001000100010001110100001000001100010001110000011101001101010000110100001110000101010000001100001011000111010001011000100110001111100010000100000110000001000000011000101101001111010011101000111001000110100010100000111110001100010001011000000011001001110011011000000000001100110001000100011000001101010001110000101101000011010000101000011100000010000000101000010001000011100010111000100100001100110001100100100100000011100010110000011001000001000000110100100011000100010010101000010010001010010011001000110101001101010000010100001100001000100011001100000000000101010000101100001001001101110001001100110100001001100001100000101100001001000001100100000101001001010011011100010111001110110010011000110001000100100011011000101011000001100000110000100100000111110010000000100001001100010001111100011000000010100001110000110010000101100010010000000010000111010010101000011101001100100000011100000001000011000011000000000110000111000001000000010110001100010001011100010000000000010011010000010111001011110000000000100000001110110010010100011000001000000000111000000000001000110001111000100111000000100011001000010110001110010000000100011100000011110010101100010010000011100000000100011100000111100011011000001100001010010001011100110010001100000001010100100010001101110000101100001000000011100001100100110111001101110011011000001010001100010000010000000001000111000001100000100110001001100011110000001010001100100000011000110111001001000001000100100011000111000001101100011101001100110001000000001101001110110000001100111011000101110011010100111000001111000000111100010001001000000011101100110111000011010000000000011110000111110010101000000001001000000001001000101010001001110000010100011100001110100010110100011000000000000011110100000011000010110001010000110011001001100010000100100110001101010000101000111000001100010000110000011010000010010001111100110011001011100010110100001011000110010000111000110010000010000011000100101000000111010011101000010100001101100001101000011111000111000001110100101001001100100001000000110111001001100010010000101000001000010011011100111000001100000010100100100110001011110011000000010111001010000011011100001111001100100000001100110011001010100000010000000101001111010000000000011111000101000000000100111010001011100011110000110111001011110001111000000110001011010010101100000111000111000010000100101111001101100001100100101001000000110000000100000000000111100001101000000110000000000001001100110011001101010001001100010110000110010001110100011101000101110010111000000101000011110000011100110101000011100010100000101000000010100000011100011110001101100010001000100101000000100011010000101001000001010010001100101100001000100010010000110001001010100000100000001110000111110000101100001001001110010010010000001100001011100001101100100010001001010010111000110111000000000011001000101010001110110010000100100000001110110011011100011111001110010011111000010110001110000011100100000001001101010001000100110110000110000001000000100100001111010010000000010011000001110011011000010110000111100001011000111001001010010011000000111011000100000001110100010011001000110000110100100100000101100010111100101111000110100010011100000101000111110010110100100100001001110010101000111111000101100001111000011000001101010000010100100011000110110010000100111111001100100011000000010000000001110011010000110010001101110001111100000001000111100010100000010001000110010000001000110100001100110001111100100000001100010010110000100010000100110000101100011101001011110010010100111000001001010000100000000100000001110011101100011100001011000000101000111000000111000010110000001100000000100011010000011011000100100010000000110000001011010000101000100111000100000010101000001110000110010011111100100100001000100000100100111010000110000011000100111000001101010000100000011010000110000011010100101110000000000010100100010111000011000010001100111101000110100011111100100101000001100000001100001101000100100011100100101000000010010001101000001101000111110011001100101110001100010000011100111010000111110011100100001001000010110011000100101111001110110001011000011101001011110010110100110110001101100010011000010111000110010001001000100100000000110011100000100000000010000010011000100001001010110001000000111001001011110010011000010111001101110010100100100110001110010000010100111111001101110010111100111110001100010001100000000010001011010001100000111001001011010001110100111101000110100010111000101001001001110011000000001000001110000000111100100001000110100010100000000001000101010010110000011101001100010001011100111000001101000001001100010101001110100010010000001001000111100001111100110000000011000011101100011000000000100000100100000110000111010011001000101101000100000010111100000000001101010000110000010010000001100001110000101001001111000000010000000100000111010001010000100111000111000001000000001110001000000000000000010001001010110001000000110101000001100011011100110110000011000001000100111110000011100001000100011000001101100010111100000110000111110011111000101000000110100011011100111010000010000010000000100111001011010000001000010101000000000001101100110110000101100011011000000000000111010010001000111111001010100000000000011100001000100001010100001010000001010010100100011101001011010001110100100110001111100001001100001001001101100000010100001010001010010000011000010100000001000010000100011101001101100010001000000100001110010001010000101010001010100001011000011111000111010010100000011100000111110010111100010011001001010001010100110011000100010011011100011100000101000000010100011000000001100011111000110111001100010000110100011010000010110011011100011011000110000000100100111111001101110010110000001010001001000001010100000101000110010011110100100010001001010000001100100101000110000000100100111101001010110010000100000010000010110011001100101001001001110000010100111100000101000001100000101101001010010010000000000000001111000011100100111100000110000000001100101001000101110010110000000000001011010010101000011100001000100000101000001010001000000000001000111011000101110011101100100001001010100010111100111111001001100011000000110100001010010001110000110001000100000010001000101001000001010001111000001101000101100001101000100110000111100001001100001100000101100011100000110110001110000011100100000110000101100001101000001110000100000011110100110011001001010011011000100111001000110000010000000010000010110001000100101101001101010010011100010001001101000011101000011011000110000001001100100101000100010001111100011110000011100011111000001100001011110000101100101011000011100010101100000110000011100010110100000110000111110010011000011111000100110010110000010111001011100011111000010100001101100000101000111001001100110001110100011111001110000010001000111101001011000001111100100000001010000000001000001000000011000010000000001111001111010011001100010111001110100011000000101101000001100010001000000000001010100001010100010011000000100000001000101000000010010011111100111111001101110000111100110100001010110000100100111100001100100010001100011000001000010010001100111101001110110010000100111000000010000011010000000111001010110010100000111110000010110000001000100011001101010000010000110101000111000000101000100001001001110010010100010010001110000011101000010101001101110010100100000011001010110011100100100100001000010000000000110101001010100011101100110111001001010001110100011111001001100001101100011110001000000010101100111111001010110000011100011010000110010001001100110101000010010001000000101001001110100001011000111000001111000000111000010100000111110001111100100101001010010011000100110000000000010010110000110001001000000010010100000000001101000001010000001111000100010011101100111100001111100000111000100101001111000001010000011110000010110010101000100011000100010000010000001110001101100010001000011101001101100001011000111011001100100001110000100001000001010000001000001110001110010010111100001110000111100000000000001001001011100011110000010110001000000000010100001111000111000011101000100001001000010000000100100011000010010001000000011000000101000001111100010100001101110001000000101010001010110000000000110100000110100011001100101001000100100001001100001100001001110000010000110110000110000010011000111000000100010010010100011101001001010000100000000101001000100011100100010000000111100010001100101011001001110010010000101110001110010001011100011011000111110011011100101110000100010010000100111001001000110000111100011110001000100000010100100001000101110000101000110001001000100000101000010100001010110010110000111011001011010001010100100010000001000011100000000001000011110000101000100111000100110000000000001000001100100010010100100011001000100000011100110011001101010000101000001111000110110001011000111011001101110010111100001000000100000000111100111111000000110011001100111001001011010000010100100111000011100010010100011110000011000001100000101011001100100011000000000100000100010001111000010000001110100010110000101011001010000011000000001101001110010000110000000011000100010000100100100100000110010011010100111010001001110010111000101100000011110001010100001110000101110001000100110010000101100000101100110010000110000011110000101011000011010000101000001010001000010010010000110101001001110010110000100101000111100001100000011101000111100001010100001011000101100011010000111011000000110001010100001001001100100011111000001110000000110001111100110001001110010000010000010101001110100011100000001100001101010000101000001110000001110000001100101101001110110011111100110010001000000001111100001011000100000010110100111100001100100010001100011110001111000000110100010110001111110010001000000001001101010001100100110010000111000000011000011110000011000000001100110010001010010010011100001010000000100011011100101011000101010010110100111110001011010011111000100110000000100010011000001100000010100011111100101100000001010001100000011110000111000010110100100000000111010010110000100011001110110010011100111111001001100001010100110010001001100010110000110010000100100000101100110111000110110010101100011101001100110001100100000111001111110000100100110001000101000011111100100110001100010011111000001100001110110001001100001110000110110000001000000010001000110000100000110100000010110010111000101001000000010010010100100100000000010010010100000101000101000000000000100110000001110011000100000001001100100000100000001000001010000001001100111100001010110011011000111011001011010010100000011111001110010011001100111000001011000011011100111011000001000000001100111111000111100001011000010101000010100000001100100011001111010000010000110101001000010010000100111010000111000000110000110101000100010000100100010101000010000010101000000000001111100001101000101001000111110011010000101100000110110001110100100111000111000010100000001001001010010001000100111010001101100010111100000110001010010001000100000100001100000010101000011001001011100000101000100000000010000001010100011011000001110000010000101101001010000000100100000111001000000000000100110110001010100001011000000111001001010001101000111101001110010010110000011101001110110010000100000111000011110000001100001000000110000000110100111111000000000011101000000001001001000000000000111011000110010001110100001010001000000000001000111010001001110000101100011110001110010011101000100000000100010011101100101101001000010011101100100010000111010000110100110000000100000000110000111011000011110000011100101110000110110011010100111010001000010011101100010001000100000011011000111011000010110010110000110111001011110010111100101001001110000000000100011110000110000011100100101000000010000010011100001101001001000010100000100101001100010000010100111000000111000010101000111011001100110010010000110001001110100010000100001011001010110011110000001001000001010001101000100111000011100000101000111011001100100000001100010011001111000011000000010110000000100010100100010010000001000000111100111011001111010000000000000001001010110010101100110101001000010011001000101101000111110011000100001001000000010010111000011011000011110011100000011001000111110011110100001001000010110011110000100001001010000001010000101111000101110000010100100001001000000001011000000110000111010000011000011001001000010011101100110110001111010010010100110111000100010000111100011011001010100011100100011101001101100011101000000100001110000011100100111101001111010000100100000100000010110001011000100110001011010001011100100100000000110010011100111000001000100010100000110111001010010000111000110101001010010011001100100010000001110001001100011001001111010010010100000010001100000000011100010010000110100001100100011110000100010000000100111110000001100011010100110101001101000010000000001011001011110011010100010010001011110011001100010000001111010011010000001001001010110000110000000111001110110001100100100001001100110011111000000001001000110001010000101000001010010000101100110000001111100000101000111001001111000011011100100001000110110000001100101011000110000010000000100001000110010000101000111001000011000001011000010110001101110001101100011001000011000010101000010100001011000001110100100001000010010010101000001000000001110010000100000110000111100000001100001111000001010001101100011101001001100001110100100100001101000000110000011111000001110001011000001110000000000000101000011011001100000011010100000101001001110010010100111010000111010001010100001101001011010001011100000110001010000000001000100000001000110001010000001110000111000000111100001111001001010010001100111000000000000001100100101110000111110001000000010100001010010010011000110110000100000010111100010100001011100010000000111111000110100010110000101111000110000001110100110101001111100001001000010011000000000001011000101011001100100001011000011000000011110001000000100101000001000000000000100010001100010001000000101001001101010011011000111001001100100000111100000110000100100001110100001101001011000011100000001100000110100011011100000100001001100011110000010011000010010010011100000000001000110011000100000011000010110010011000001011000101000000101100001100000001100010011100000100001010000001111000100010000000010010011100111001000100100011101100000010000000110000001100111010000111010001110000000000001011010000111000100001000000100010011000111001001101110001010100110111001001000011000100100011001000100011011100101101001011000010100100011001000000000011101000111010001111000001111000101000001110100011011000101110000111010000010100100000000010000011100100000111000001110001011100001001001000010001100100101000001100000011010100000010000110110011010100010100001011110010011000100101000011110000001000100101;
		
		// Wait for global reset to finish
		#100;
				
		// Generate a reset
		CPU_RESETN = 0;	#20;
		CPU_RESETN = 1;	#20;
		
		BTNC = 0; #20;
		BTNC = 1; #20;
		BTNC = 0; #20;
		
		// Give a long time for machine to finish
		//#8000;
		//32000;
		#500000;
		
		// Wait for global reset to finish
		#100;

	end
		  
endmodule

