`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   20:12:24 10/05/2015
// Design Name:   quickhull.v
// 
////////////////////////////////////////////////////////////////////////////////

module quickhull;

	// Inputs
	reg CLK100MHZ;
	reg CPU_RESETN;
	reg [4095:0] points;
	reg [7:0] SS;

	// Outputs
	wire [4095:0] convexPoints;
	wire [7:0] convexSetSize;

	// File
	integer file_results;

	// Parameters
	parameter CLK_PERIOD = 20;

	// Instantiate the Unit Under Test (UUT)
	quickhull UUT(
		//Inputs
		.CLK100MHZ(CLK100MHZ),
		.CPU_RESETN(CPU_RESETN),
		.SS(SS),
		.points(points),
		//Outputs
		.convexPoints(convexPoints),
		.convexSetSize(convexSetSize)
	);


	initial begin : CLOCK_GENERATOR
		CLK100MHZ = 0;
		
		forever begin
			# (CLK_PERIOD / 2) CLK100MHZ = ~CLK100MHZ;
		end
	end	
		
	initial begin : STIMULUS
		
		file_results = $fopen("output_results.txt", "w");

		// Initialize Inputs
		// === Small input: 15 points ===
		CLK100MHZ = 0;
		SS = 15;
		CPU_RESETN = 1;
		points = 4096'b0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000000000000000000000000000000000000000000000000000
					   0000000000000000
					   0000011000000110
					   0000010100001000
					   0000001100000111
					   0000011100001001
					   0000011100000100
					   0000001000000101
					   0000010100000001
					   0000010000000110
					   0000010100000011
					   0000010000000010
					   0000010000000101
					   0000010100000110
					   0000001100000100
					   0000110000001001
					   0000101100000001;

		$fwrite(file_results, "Points:     ");
		$write(file_results, "Points:     ");
		integer counter;
		for (counter = 0; counter < convexSetSize; counter = counter + 1) begin
			$fwrite(file_results, " %h", convexPoints[(16*counter)-1 : (16*counter)]);
			$write(file_results, " %h", convexPoints[(16*counter)-1 : (16*counter)]);
		end


		// Wait for global reset to finish
		#100;
				
		// Generate a reset
		CPU_RESETN = 0;	#20;
		CPU_RESETN = 1;	#20;
		
		// Give a long time for machine to finish
		#5000;

		// === Medium input: 50 points ===
		//Input next test
		SS = 50;
		points =  4096'b0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						0000000000000000000000000000000000000000000000000000000000000000
						00000000000000000000000000000000
						1001101101010010111001110111011001101100100000101010001001001000
						1101100111110010111010110011010000000100001011110000001011110010
						0010011100100100101101011100101111000011011011010001100100111011
						1000110000001111100001111101011010011101010000011011011011011101
						0110010111011010011101010100001110101101101001110101101010101011
						1111001000111000101001011111100111111010001101000010100110101011
						1000111001110111011010000100001010111100010100100010110001110000
						0000010101011001010110101101011000100010010111001101011011110110
						0100100101010001011100011000000001011000011100100101110010000111
						1101000100110010000010001000111010101001011011101000101111101111
						0111111000111110011011001001001010001010000010101001100011100000
						1010000011000110110110001110001011100011100111010010101101010110
						01011011011010100100011110000011;

		// Give a long time for machine to finish
		#5000;

		// === Max input: 256 points ===
		// Input next test
		SS = 256;
		points =  4096'b0101110111110101111110100000100001100000111110100110001101001011
						0110100000101100011100011000000110000111110011010111011000010101
						0001010000001011100011110001100010111010111001110100010010101011
						0010100100010111100111000110011000010010000110010111111010000011
						0001000000011101111011000011100011000011100001000101101111101001
						1001101101100000010001011000100100101110000111111010010110100110
						1101000010010001011110001010100000100001010111011101110011000011
						0010000011000110011110101110001100100001011111011101101101010000
						0001101100110010011111001010110110001111101001010100100101001011
						0111011111100100100100001111110011111001100010000110100101100011
						1010100010100010110001100100000101101011100010110110010010001000
						1110001100010011001100010111101001010001010010111010001001100011
						1011011001011011011100000011010001100101110111101111111100101010
						1011010011000110101110001000101011101010101111001111000000100111
						0110101110111000010001101101101011011100010110011110000111111010
						1110000111010110111111011101010100100010011001010001111000110110
						0100111101100101100001000010000100011101001101101111010000000000
						0101101011000011110110000111101000000110011111101010111011101011
						0010110010110100110100010101000001010000011110001100101001010001
						0110111001001101110010110100001000110010000010010000111010100100
						1010001101010000111010001110000000010110111100011000011000000100
						0100100110000010010001100101000011001111011010110010111010100110
						1111010001010001111011110010100100111011001101110100101111100011
						1101101000000001001111111010001010001001001101011101010110111000
						0100000010110000111000110111000011111000001011001101100010110110
						1001010101001110101101000000110100001001001101001010011001000101
						1010100001001011001111110001101111000100110100111000111000011001
						1000001101001010011011011110000000100001001010100010001101100101
						1110111100110011110011110010111100111101010010010110110110111110
						1111000010011001111010110101011101001110111001101110101011110111
						0010111101110101110010011110001000000111010010100001110001001001
						0100010101001100011101100010110100011101111100110001001110001101
						1100111110010011111000010000011100010111011011101111010110000100
						0001011111000100001100000111010110000010010011011101100100111000
						0010110111000110101111110010110101011010000111100001111000010010
						1001000111111001100111101111101100101011111111111011110110100010
						0111110101011111111001000111110011000111110110000000101011010111
						1010101011011010001111101000000000011011111001101011100110100010
						0011101001010111010110100101000001111011110100011100001100000111
						0101100010100110001001000000100001010000010101110011011001110110
						0110101001100010010000010011010101011110111101110110110111111110
						1011010001110101100000001101001000101110000000000010010100001110
						1001010000000001110001101111100001000010100100001010111001010100
						0101011001001010011110100100000000100111110000101010111010011110
						1001101011011010001010101010011101111100100010100001011010011100
						0010000001010001011001011000100011111001010010000011100010001011
						0010011000001101000010110001101000110011010001101100000010011010
						0010111111111101101010110010111011101011101000111000110100101111
						0010111001000101100010000011101011110011001001100110011100001010
						0001111000110011100011011010100111101000001000111000011011111010
						1010111111010010111110000111000010100000100111111001001010100000
						0001010001001011111000011001110110010101001011000101101011100101
						1101101110011100101100110001010000110010001100100010111101010001
						0011000111011001111100100011101011111000100001010111111101001111
						1011111111010110001010000100011001101000011000111000110010010001
						1001010111000011001000100111111000001111011100111011011000000001
						1011010000101011111101000101111001100010100101110000110000111100
						1010010010001011000001000100101010011100010001101010001110001110
						0000010100001001110111001111001001101011010011011111110100011101
						0010010000110110101011111000001001101001010101010001010101101011
						1101010001100011001001111011010111110011110011110001110100110100
						0010101110110001110110011011101001011111000011001000110010101111
						0111100000100100001011010101010111001100001110111000100011001110
						0110001110101011110000001001100101100101010101011111110101011010;

		// Give a long time for machine to finish
		#5000;

	$fclose (file_results);	 

	end
		  
endmodule

