`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   20:12:24 10/05/2015
// Design Name:   quickhull.v
// 
////////////////////////////////////////////////////////////////////////////////

module m_port_ultra_tb;

	// Inputs
	reg CLK100MHZ;
	reg CPU_RESETN;
	reg BTNC;
	reg [16383:0] convexCloud;

	// Outputs
	wire [4095:0] convexHull1;
	wire [4095:0] convexHull2;
	wire [4095:0] convexHull3;
	wire [4095:0] convexHull4;
	wire [8:0] convexHullSize1;
	wire [8:0] convexHullSize2;
	wire [8:0] convexHullSize3;
	wire [8:0] convexHullSize4;
	wire processorDone1;
	wire processorDone2;
	wire processorDone3;
	wire processorDone4;
	wire QINIT, QPULSE, QDIVIDE, QCONVEX_HULL, QDISPLAY;

	// Parameters
	parameter CLK_PERIOD = 20;

	// Instantiate the Unit Under Test (UUT)
	m_port_ultra UUT(
		.clk (CLK100MHZ),
		.reset_n (CPU_RESETN),
		.ack (BTNC),
		.convexCloud (convexCloud),
		.convexHull1 (convexHull1),
		.convexHull2 (convexHull2),
		.convexHull3 (convexHull3),
		.convexHull4 (convexHull4),
		.convexHullSize1 (convexHullSize1),
		.convexHullSize2 (convexHullSize2),
		.convexHullSize3 (convexHullSize3),
		.convexHullSize4 (convexHullSize4),
		.processorDone1 (processorDone1),
		.processorDone2 (processorDone2),
		.processorDone3 (processorDone3),
		.processorDone4 (processorDone4),
		.QINIT (QINIT),
		.QPULSE (QPULSE),
		.QDIVIDE (QDIVIDE),
		.QCONVEX_HULL (QCONVEX_HULL),
		.QDISPLAY (QDISPLAY)
	);


	initial begin : CLOCK_GENERATOR
		CLK100MHZ = 0;
		
		forever begin
			# (CLK_PERIOD / 2) CLK100MHZ = ~CLK100MHZ;
		end
	end	
		
	integer counter;
	
	initial begin : STIMULUS
		
		// 16 size, 32 range
		//points = 16384'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100011000000111010001000100001100000010100000001100000000000101110000110000001001000111010001001100001000000100100000110100010011000011010001000100011111000111010001111000001000000100000000101100000111000001100000010100001001000110000000011100011001;
		
		// 32 size, 32 range
		//points = 16384'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000100001110000001011000111010001100100011011000100000000101100000010000010100000111100011111000101010001111100011111000110010001101100001010000100010000011100011010000011000000001000001100000111000000111000000111000110000000101000011000000101010000111000000110000101010001110000010101000111110001011000000101000011110000111000000011000000000000011000001101000110100001100100011111000010110000101000001010000001010001100000001000000100110000000100010011000010100001100000001001000001000001101000000011;
		
		// 64 size, 32 range
		//points = 16384'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000101000100000000110000000110000001100001010100001001000100010001010100010110000010010000100100010110000001010001111000001110000100100000111000001011000000000000011100001001000001100001100000011000000111110001111100011110000101000001010100010110000011010001000000011100000010100001101000000001000100010001100100000100000010100000111100011001000010110001001000010101000110000000101000010111000100010000101100011110000011010001001100011001000010100000000100001101000111110001110100011011000001000001111100000100000101110000011100010110000000010000001000001110000000100000011000001101000101100001101100010110000110010000110100001100000111010001111000011101000001000001101000010000000100010000110000000010000000100000010100010101000111110001011000000000000111110001000000000000000100100000100100001111000110010000010000011010000110000001110000010001000111010001101100011000000110000000110100010110000010010001100100000111000100000000000100010001000011110000011100001010000010010001111100000101000000010000010100000000;

		// 256, 32
		//points = 16384'b0001011000001111000011110000011100011000000101010000110100011001000001000000101100010111000111000001011000000011000100100001000000010100000000000000011000011101000010100000010000001101000101110001100100001110000001110000000100001100000001110000011000010010000111110000000100000100000110100000110000010111000100100001000100001010000001100000001100000011000100100000010000011101000000110000101000000100000110100000011000010000000001110000000000010011000001110000110000010111000000000001110000011100000101100000000000000101000100110000011100011110000000000000000000001110000000010001100100010001000111010001010000000111000010010000111100010110000100100001010100011111000100100001000000010100000011100000011000000011000010100001100100011110000011100001111000011001000000110001110000001010000001010000111100011000000010110001110100010101000011110000001100011111000110000001111000011111000001100000100100010110000100110001101000011101000011000001011000011001000101000000011100000011000111000001101100001001000000110001001100011100000000010001110000010001000100010000101000000100000000100001110000010100000011100000000100010010000001000000111100001100000110000000011000000010000010010000011000011111000000110001110100000101000010100000011000001011000000110000110000011110000011010000101100000101000000000000111000011111000001000000001000001111000011010000100100000111000000110001100100010010000110110000110100001000000000110000000000000000000001110000010000010001000111010001110100010000000101100000110100010011000111110000011100001010000011110001010000010001000001000000101100000101000001010001111100000010000100000000010000011111000101010000100100010011000000010000000100001011000001110000111000001101000001010000001000001100000010110001010000000110000011010000100100011110000100000001101000011110000100100000000000000101000011110000011100011010000010100000100100010000000111000001101100000010000101010001010000011110000110000001111100001011000100000000001100010111000000110001010000010010000001010001000000000100000001000001010100001101000111000000010000001101000110010000100100010010000010100000100100000000000111000000001100001100000100000001001000000101000101000000010000010010000111010000011000010111000010000001010000001111000001010000111100011100000001100000001100011011000100010001101000010100000011100000011000010011000101100000011000001100000000000001000100011001000000100000110000011011000011010000111100001110000011000001001100011100000010110001110000001001000100010001110000000111000101010000001000010110000111010001000100011010000010110001110100011110000111100001100000010111000011110000111100000111000000000001000100001001000110100000100000001110000100100000011100000110000010000001000100010100000101110001011000010100000011010001000000000001000010000001011000000101000010110001011100010011000100000000011000001111000101010000011100001101000101000000010100000100000000100001000100001010000011000000111000000110000111000000001000000010000010110000010100001100000100100000011000001101000010010000111100001011000111000000100100011010000101010001011100001011000100100001100100000101000111110000110100001100000110000001111000001111000000000000000100001101000110100000011000011100000101100001101100000110000100100001100000000101000101110000101000001100000110000000011100001001000010010000011100011110000101110000000000000000000100000000001000010101000111010000111000000010000101010001111000001001000111100000111000011101000001100000110000011110000001100001010100010111000110110000000000001001000001110001000100001100000101010000010000001000000011100000011000010010000111100001111000000001000010110000110100010110000100110000011100010101000001010001001100001010000011000001111000001100000001010000110000000001000011010000001100011110000101100000010000001001000101010001010100011111000101100000000000011101000110110000101000001111000100010001111000000000000111010001110100011000000111010001111100010001000101100000010000001010000100110001110000000111000010000000110000010100000100010000100100000001000001100001110000000001000000010001110000000001000100100001111000011000000110010001111100011001;
		
		// 16, 64
		//points = 16384'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010001111000000001000000010000100100011000100111110000000010011111000110011000000110000100000101100000100000010010100000010000100000000010000000011000010010010110000001101000011100010110100000110001111110010000000111011000000010000001100010100001011110001000100111100000100100011100000100011000011110000110100111101001001010001111000100011001001100011110100011010001111110010111000010110000111010010101000000001000110110001010100111000000100110010110100000101000001010010100000010000001101000001000100111100;
		
		// 32, 64
		//points = 16384'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010001001010001001000110101000111000001010000101001000011110001001100111101001111000011011100000110000011100010110000011001000111010001000000101000001100000010011100011001001001010001111100100011001101110000010000011111000111110010000100110001000100010000110000010100001001110010010100111111001011100000111100110101000110010011000100110100000000100010100000001101000011110000101100011011000000010001100000001001000101000001111000111101000110110010001100010011001111000011111000000011001100000001000100011100;
		
		// 64, 64
		//points = 16384'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000010101000111000010000000010010000110100010100000001101001101100000110000110011001001000010010000100111000000100000011100101101001000000010010000011110000101100011010100001000000100110001101000001110000001010000101000101101000011010010110000110101001110100000011100100111001000010010101100000000000011100011011000101010000101010001000000101111001101010011111000010100001011010001011000010100000100010011010000000111000100110001010100001001001110000011110000101001001100110000101100100101000000100001001100011111001111100000000000011011001111110011111100100111000110010001010000100101001101110001111100111100001011110011000000111100000000110000001000111111001111100000001000111111001110100010111100110100000011010000110100000110001110010011010100101011000010000010010000111100000001010001100100111011000110100011000100000110000101100000011100100110000010000001111000011001001010000001010000011000001100100000110100011000001111000010000100011100001100010010100100001111001010010011011100111110001010000000100100100010;
		
		// 256, 64
		convexCloud = 16384'b0000010000000010000011010010101100001101001111110001001000101000001100010000000100001100001011000000110100000111001001100001111100010110000010100010010100011011001010100001010000111000001010000010100100001101001001000000101100110101001011010000000100101111000001110001011000111010000101000011010000000010001011000011011100111011001100110000011000101000000100110010111000100101001110100000000100111011001100010011110100100000000000100010000100111011001100000000010100101111001000010010110100001110000110100010101100111001000110000001000000111100001111000010100100000011001011110000001000110111000000100000110100101110000011010010110100111011000100010000110100111001001001100000001000111101000111110001100100111000001001100011100100110010001001110000010100111001000010010011101100000110000001010011101100100011000100100001011100101010000010110000011100001010001111000011011000000100000100000000111100000101000110100001100000110100000110100001100000110010001010010011101000001010000010000001010000010101000000010001000100110010000110100001000000000100000110010011110100101100001111100011010100010011000000000010010000011110000110000011001000100011001011100010100100111001000011000000001100010101000110100000001100110011001101000010110100110011001101010000001000110010000100110001101000000000001111010010010000111101000111000010011100011011001101000010011100011100000101010000111000001000001110000001001000011100001100000001111000011010000100000000100000111100001100000001011100001111001011100001001100110100001110000011111000011111000100100000000100011011001101000010010100101010000001000000011100011000000011000000001100111000000011010000110100001110000010100010101100110111001100110001110000110101001010110011001000010011001100100001000000111001001111010000010100101010000111110010100100111100001011000001101000001100000100010000110100111110000110110011010100110110000000100010000100101100000000110010001000100101001000010010011000110110001010100011101000101000001101010011000100000011001000010011100000111001001000010000101100111010000101010001110100101111001101100000101100010100001110000000100000111000001000100010111000010011001110110001100100100111001011100010001000000100000111110001100100000101000111010011001100011101001010110010110100001110000101010000011000011011001110000010011000011000001000010011010000100101000110100011111000010110000000100011110100011011001001110000010000100111001111010000111100011000001010000001110100011101001111010000000000011110001010010010100100001100000001010001111100101100000110110000100000101101000000010001001000001101001100000000000000100000001111000001100000111010000011000011000100100001000101010001000000010000001101000011100000010100000011000000010000111111001010000000100100000101000110100001000100001100000111010001011100000000000000110000100100000110000111110010011100011011001001000001001100011110000010000000110100111110001000110010010100011000001000100011110100000011001101000011101000110011001011000001001000110011000000000011111000000100000111000001000000010110001100010010000100001011000010110010111000111101000111110001110000010011001000000001011100001100001100010000101000000001001110010000110000011111000001100000010100010111001011100001110100101111000010100010111100001001000011000011010000000000000001010000000000111001000011000000110000011001000000100001010100110110000101110010000000010000000111110000001100110101000001010011000000100101000111110000010000100101000101100010010100000100000000100010101000001101000001100001011000111001000101010011011100000100001001010011110000111001001011000000000100100111000011010001101100011000000001100000101100000100001011000011001100111110001011010011001100000111000110010000000000100111000010110010111100110010000100000011011100000000000011000001111100100110001101000010110100011100000100000010101000101110001110000000101000000000000010010001111100011010001000010010001000101011000010010001100100011111001010010001000100011111001000000010000000100000001111000010111000101100000010100011101100011010001000100011010000100001001100110010010000011001000010010000010100110010001010110010011100011100000101010010110100011100000101100011101100001001001011000010000100000101001011000011110000101111001010000011101100000001001001110000001100111000001010110001111000101011001100110010010000010010001110010001111000110101001011000001010100100001001000010001111100010000000001010010000000000011000000110001101100101000000010110000100000111101000001000010101000010010000110100011110100101000000011100011110100011100000010000000000000111101001111110000100100101110001111110001110000101101000111010010101100001011001010110001100100011001000000110001000000011111001110010011111100011111000101100000111000101101000100010011100000100100000101010000111000011011000011000011111000000000000110110011011100001000000000110010010000010010000110010011010100010000001111000000100000111010000100000010111000001001001100000010111000111011000000000001011000000010000010000011010000101000000101010011000100100001000100000001001000000111000000110001111000010011000000110011001000111110001000110000000100111100001001100011100100100001000000100001001000001101001110110001100000010000001011010000101000010010001100110000000000010001001001100001101000110111000110010010010000101000000010110001010100111000000111110011101000111100001110010010010000010101001111000001000000100100000011010011001000000000000100010010100000010011000001000000100100100100000101100001001100101100000100010010110100101000000101000001011100000010001010100011001000111111000100110000111000111001000000100000110000110010000101110000001000110100000111110010000000110101001110000010111000001111000101110010100000111000000100000001101100010001000101110000000000010011001100110010000000000100000100000000001100110110001111100011010000001111001111000011001000010010001011000011111100010001001000010000000000001011000000000001010100110100001000100000100100011110000000010010011100001110000000010001111100000101001101100010001000111000000101110000100000100011000110110000000100110111001101010000111100101011001000110001010000100111001010010000010000000010000101110011011100100101001010010001100100111110000001010000101000110001001010100010000100111011001010110010111000111010000111000001111000010101000111010010011100001101000111110010000000010111001011000010111000111101000100100010110000011001000011110010001000010011001110110011001100011001001101010011100000110001001000000010000000100011001100110001110000010100000000110001010100011011001111000000011000011110001111010011110100110000000011100001101000110111001000100000011100101110001001100011010000101010001100000010110100100010000001000010010000001110001110010010100100010101001011110011110000011010001110010000011000101110001111110011101000100111001011110011000100011001000011010010111100111111001001100001010100011110001010100000001100110110000100000011001000110110001100110000000100110000000110110000111000101100000010110011110100100101001100100010010100000111000110100000100000001111000001000011011100011100000001100001100100010010001101110011000100010000000100000010001100001001000110110000111100000111000001110000010000101100000100110000110000100110001001000010001100110100001111110000111000000001000001100000111000010010001000010010100100011101001101110011010000010101001000000010010100001011000100000001011100001110001110100010000100111111000100010001010100111000000000000001010100111110001101100010011000001010001001100010011000111100001010000011010100001100001101110011101100111011001011100001000100010100000111110010101100000010000111010000101100101001001011110010000000001000001000000000001100001010000100100000011100010101001110010000101000110011000110110001000000100010001100110000110100000110001100010001011100110101001001010001111100101100001010010001001100110101001001100011101000100001000101010010111100111000000011100010001000110011001010100011111100101101001011010010101100110101001001010011111000100101000111100010001100011111000000010001100100000000001110000011101100110001000101010000000000000100000001000010110100010000001010000010110000000100001100000010001000011000000011110000110100010101001001000010101100001000000111000011110000001111001101000001010100111101001011000010111000100010000010010010001100101101001010100011010100010010000001000011100000100110001100110010100100110011001001000000000100110111000010000000001000111111000110000001110100001100001101110010111000110001001110000011101000011111001000000001110100011101000000010001111100110111001110100011111000101010000100100001010000011011000010110000101000010111000111110001101100111011001001100000001100000000000101110000000100100000001100110001110100010011001100010011110000010000001111000001001100101000000100000000000100100011000011100000000100001001001001100011100000001001001011010010100100001000000011010010010100011001000110110000000000011101000001100001101100010001000000000011010100010010000001100000100100011001000010000000001000111010001101000011101100011000001110010010001100001101001110100000010100011011000100010001001100011100001001010010000100010111001010110000001000110110001011100011000000110101000010100011000000100100000101000001111000000101001010110010111000001010000101110011100000001111001010100000111100011010001101100010101000111111000110000010010100001100000111010010000000001001001010100010111100010011000111100011010000111010001100100001011000011111000110000011101000001001000100110010100100000011000101000011111100100000000101110011001000011001001111110010111100100000000100000001000000011010001110000011100100110000001011000011100100000100001001010010110100000101001010100001010000011011000001110010010000111100001110010010101100100101000001110011111000101110000101010001110100110001001011100000000000000101000100000010111100111011001011010000111100100111001100100011101000101111001110010011111100010010000100000000111100000000001011010001110000011111001001000000101000000100000111100010110000001101001111000000010000010101001101110001000000010110001010010000110000000111000101000011101100101110001000010000010000110011000111010000000100010001000011000001010100001110000100110011110100100110001010000001000000001111000010110010101000011110000110110000110000000100000110000001100000000110000011110011010100001110001011010001111100000111000001000010110000011010001110110000111100000111000001000010010100100010001101100011010000000100001001100001011100110011001101010010100100100110000101010001110000100111000000000010010100100100001100110000000000110010001010000000010100100110001101110010101000111000000100010001001000101111000110100011101100000110001000010010111100011111000111000001001000010000000000000001001100010100001100110001101000101100001111100001111000110101000011000000101000011000001001110011100100000010001010110000110000001011001000100001111100110010000011100000000000000101001011110010101000111000000001110000011000101101001101100001100000011100000010010001100000101011000000000001110000001111001110010000001100001010001000010000111000110000001110010001000000011110000100000010000100010010001001100010010000000100001100000000001000111011000001110011100000011101001111000001001100101101001100110010010000001101000100000010010100101101001111100001110000100001000101110000001100111010000010100001010000110110001101000010000100011100000101100000101100111011000100100011001100101000001010110000110100111100001100100010111000000001000011110001010100100001000110100001000100001011001110100001110000110110001100100010111000001110001101100000110000100001001000110011000100111111000100100010000100010110001111010001101100100101001110010001110100001111000011100010101000001101001110110001001100010100000101100000010100011100001001010001001100010010001110000011000000001101001110010000100100111000000000000010010000010000000000100011001000011011001100110001101000100101001100110000000100100001001010010011100100110011000011000010100000010010000101010001001000100011001010110000010100001000001110000011001100111010001111000011000100011100001111110000011000111001001111110000010100011010000100110000100000110111001110000010100100111011001111010000101000011110001000110000011000110110001110000000100000111100000000000001101000100110001110010001001000010100000111010000100000001111000110110000111000111010001101110000010000100011001010000010111000011011000000100000000000100000000011100011110100110001000111100001100000110000001100100011001000000101000001110011111000111000001100110010001100011000001101010000000000100000001110100010000100100001000001100011111000000101001101000011011000001100000110010010100100011001001001110001111100101110001010000011110100011010001111110011010100101001000101010011101000100010001110000010100100001000001101010000001000000011001100100000001000001110001001000000101100111001000000110000011100011010001100010011110000100101000110010010010000010110000010000010011100010010001100000000101100000101001100100000000000101110001001010001011000011100000000000011111000011100001111100010100000110000001011100010110000001001001011010010100100010011001110100000001100001110001000100000100100011010001101110011100000011110001100010011101000100100000011110011000100110101000110000000000100010100001111110011001000100011001011100000001000001010001010100010001100001000000101100010100000101011000010110001100100001110001111110000100100111001000000100011111100111011000101110001000000100100001000100001010000100000000010100011110000010000001000100011101100101101001000110010000000010100001100110001100000001110000100110011100100110000001100000000110000101111000101110000101000111111001010110000101100001110000010010010100100011010000100100000011100001100000111100000111100111001000111110000000100010000001000110001111000001100001100100011100000011110000111100011010000101001000100000001001000001100001001100000100000101000000111000000000100110010000101000011111000111110001101000011001100011101001110110001011100100011001010100001000100001001000000010000001100101100001110000000001000000111000101110010111100100001000000010001010000100110000001010010000100000011001011010011000000010101001010010011111000001010001010010000000000010101000010010000100000100111001011110010011100111010000001000000000100000010000101100010011000001111001100100001111000100110001100000001001100001100001100000000001000100000001011100001001000110000000111010010011100010000001011110010110100011111000101010001100000000000000000010001011000011101000001000011111100001000000010110010000000100110001111110001101000100001000110010001100100000111001100010000001000000100001011110011000000010100000011010011101000010011001110110011111000010011000001010000001000011101000100010010110000011001000011010000010000010000001011100001101100101000001010110011000000001111001011100001110000101111001110110010001000001001001100110011010000100001000111000010101100110100000100010000011000010000001001000010011000101100001110100011101000010111000001110011000000111110000001010000111000111101000010100000001000110010001100000001100000110010001110110000110100110100001000110001110100010011001100110010110100010111001010100010000000111001000101000000101100110110001101010000100100100000000110110000001000100000001000010011011100110100000001100011100000111000001000100000001100111100000111010010110100010111001010110010101100110001001110010001110000011110001000010011101100110001000001010011100100001011000111000010111000000101001101010010100000000010001110100010101100101001001010100010001100100110001111000011001100000001001100010011111000111101000011100001010000101011001100110001011000111011001001100001010000011001000111100000111100011001000111000010101100101111000001110011000100110100001110110010111100110101001001100001111100110010000101110011011100100000001011100010101100101111001111110001100000111111000111010001000000101101001110110000110100000101000010110010100100110001001000000000101000110010001101010001101100001001000111010011111000000111001000100010111000110100001001110001110000101001001000100001010000100111001010000011000000011000000010010010100000101101000111000011000100111000001000000001101100001110001001100011001000010011001111110011100100010010000011000001001100110100001001010011010100101001000100000011000100110100000100100010001100101000001000110011011000101110000010100001110000011110001110100000010100010010000101100001011100001001000110110000011000101010000011100001011100011001000101110001000100100100000100010000111100111000001010100010010000010010000000010010111100100001;
		
		// Wait for global reset to finish
		#100;
				
		// Generate a reset
		CPU_RESETN = 0;	#20;
		CPU_RESETN = 1;	#20;
		
		BTNC = 0; #20;
		BTNC = 1; #20;
		BTNC = 0; #20;
		
		// Give a long time for machine to finish
		//#8000;
		//32000;
		#500000;
		
		// Wait for global reset to finish
		#100;

	end
		  
endmodule

