`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   20:12:24 10/05/2015
// Design Name:   quickhull.v
// 
////////////////////////////////////////////////////////////////////////////////

module m_quickhull_tb;

	// Inputs
	reg CLK100MHZ;
	reg CPU_RESETN;
	reg [4095:0] points;
	reg [8:0] SS;

	// Outputs
	wire [4095:0] convexPoints;
	wire [7:0] convexSetSize;
	wire [8:0] positiveCrossCount;
	wire [31:0] crossValue;
	wire [15:0] lnIndex;
	wire [8:0] ptCount;
	wire [31:0] currLine;
	wire [15:0] currPoint;
	wire [15:0] furthest;
	wire [15:0] xMinPoint;
	wire [15:0] xMaxPoint;
	wire signed [31:0] furthestCrossValue;

	wire QINITIAL, QFIND_MAX, QFIND_MIN, QHULL_START, QCROSS, QHULL_RECURSE, QEND;
	// File
	integer file_results;

	// Parameters
	parameter CLK_PERIOD = 20;

	// Instantiate the Unit Under Test (UUT)
	m_port_ultra_quickhull_processor UUT(
		//Inputs
		.CLK100MHZ(CLK100MHZ),
		.CPU_RESETN(CPU_RESETN),
		.SS(SS),
		.points(points),
		//Outputs
		.convexPoints(convexPoints),
		.convexSetSizeOutput(convexSetSize),
		.positiveCrossCountOutput(positiveCrossCount),
		.crossValueOutput(crossValue),
		.lnIndexOutput(lnIndex),
		.ptCountOutput(ptCount),
		.currentLineOutput(currLine),
		.currentPointOutput(currPoint),
		.furthestOutput(furthest),
		.furthestCrossValueOutput(furthestCrossValue),
		.xMinPointOutput(xMinPoint),
		.xMaxPointOutput(xMaxPoint),
		.QINITIAL(QINITIAL),
		.QFIND_MAX(QFIND_MAX),
		.QFIND_MIN(QFIND_MIN),
		.QHULL_START(QHULL_START),
		.QCROSS(QCROSS),
		.QHULL_RECURSE(QHULL_RECURSE),
		.QEND(QEND)
	);


	initial begin : CLOCK_GENERATOR
		CLK100MHZ = 0;
		
		forever begin
			# (CLK_PERIOD / 2) CLK100MHZ = ~CLK100MHZ;
		end
	end	
		
	integer counter;
	
	initial begin : STIMULUS
		
		//SS = 16;
		//SS = 32;
		//SS = 64;
		SS = 256;
		
		// 16 size, 32 range
		//points = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001001100011000000111010001000100001100000010100000001100000000000101110000110000001001000111010001001100001000000100100000110100010011000011010001000100011111000111010001111000001000000100000000101100000111000001100000010100001001000110000000011100011001;
		
		// 32 size, 32 range
		//points = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001000000100001110000001011000111010001100100011011000100000000101100000010000010100000111100011111000101010001111100011111000110010001101100001010000100010000011100011010000011000000001000001100000111000000111000000111000110000000101000011000000101010000111000000110000101010001110000010101000111110001011000000101000011110000111000000011000000000000011000001101000110100001100100011111000010110000101000001010000001010001100000001000000100110000000100010011000010100001100000001001000001000001101000000011;
		
		// 64 size, 32 range
		//points = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000101000100000000110000000110000001100001010100001001000100010001010100010110000010010000100100010110000001010001111000001110000100100000111000001011000000000000011100001001000001100001100000011000000111110001111100011110000101000001010100010110000011010001000000011100000010100001101000000001000100010001100100000100000010100000111100011001000010110001001000010101000110000000101000010111000100010000101100011110000011010001001100011001000010100000000100001101000111110001110100011011000001000001111100000100000101110000011100010110000000010000001000001110000000100000011000001101000101100001101100010110000110010000110100001100000111010001111000011101000001000001101000010000000100010000110000000010000000100000010100010101000111110001011000000000000111110001000000000000000100100000100100001111000110010000010000011010000110000001110000010001000111010001101100011000000110000000110100010110000010010001100100000111000100000000000100010001000011110000011100001010000010010001111100000101000000010000010100000000;

		// 256, 32
		//points = 4096'b0001011000001111000011110000011100011000000101010000110100011001000001000000101100010111000111000001011000000011000100100001000000010100000000000000011000011101000010100000010000001101000101110001100100001110000001110000000100001100000001110000011000010010000111110000000100000100000110100000110000010111000100100001000100001010000001100000001100000011000100100000010000011101000000110000101000000100000110100000011000010000000001110000000000010011000001110000110000010111000000000001110000011100000101100000000000000101000100110000011100011110000000000000000000001110000000010001100100010001000111010001010000000111000010010000111100010110000100100001010100011111000100100001000000010100000011100000011000000011000010100001100100011110000011100001111000011001000000110001110000001010000001010000111100011000000010110001110100010101000011110000001100011111000110000001111000011111000001100000100100010110000100110001101000011101000011000001011000011001000101000000011100000011000111000001101100001001000000110001001100011100000000010001110000010001000100010000101000000100000000100001110000010100000011100000000100010010000001000000111100001100000110000000011000000010000010010000011000011111000000110001110100000101000010100000011000001011000000110000110000011110000011010000101100000101000000000000111000011111000001000000001000001111000011010000100100000111000000110001100100010010000110110000110100001000000000110000000000000000000001110000010000010001000111010001110100010000000101100000110100010011000111110000011100001010000011110001010000010001000001000000101100000101000001010001111100000010000100000000010000011111000101010000100100010011000000010000000100001011000001110000111000001101000001010000001000001100000010110001010000000110000011010000100100011110000100000001101000011110000100100000000000000101000011110000011100011010000010100000100100010000000111000001101100000010000101010001010000011110000110000001111100001011000100000000001100010111000000110001010000010010000001010001000000000100000001000001010100001101000111000000010000001101000110010000100100010010000010100000100100000000000111000000001100001100000100000001001000000101000101000000010000010010000111010000011000010111000010000001010000001111000001010000111100011100000001100000001100011011000100010001101000010100000011100000011000010011000101100000011000001100000000000001000100011001000000100000110000011011000011010000111100001110000011000001001100011100000010110001110000001001000100010001110000000111000101010000001000010110000111010001000100011010000010110001110100011110000111100001100000010111000011110000111100000111000000000001000100001001000110100000100000001110000100100000011100000110000010000001000100010100000101110001011000010100000011010001000000000001000010000001011000000101000010110001011100010011000100000000011000001111000101010000011100001101000101000000010100000100000000100001000100001010000011000000111000000110000111000000001000000010000010110000010100001100000100100000011000001101000010010000111100001011000111000000100100011010000101010001011100001011000100100001100100000101000111110000110100001100000110000001111000001111000000000000000100001101000110100000011000011100000101100001101100000110000100100001100000000101000101110000101000001100000110000000011100001001000010010000011100011110000101110000000000000000000100000000001000010101000111010000111000000010000101010001111000001001000111100000111000011101000001100000110000011110000001100001010100010111000110110000000000001001000001110001000100001100000101010000010000001000000011100000011000010010000111100001111000000001000010110000110100010110000100110000011100010101000001010001001100001010000011000001111000001100000001010000110000000001000011010000001100011110000101100000010000001001000101010001010100011111000101100000000000011101000110110000101000001111000100010001111000000000000111010001110100011000000111010001111100010001000101100000010000001010000100110001110000000111000010000000110000010100000100010000100100000001000001100001110000000001000000010001110000000001000100100001111000011000000110010001111100011001;
		
		// 16, 64
		//points = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110010001111000000001000000010000100100011000100111110000000010011111000110011000000110000100000101100000100000010010100000010000100000000010000000011000010010010110000001101000011100010110100000110001111110010000000111011000000010000001100010100001011110001000100111100000100100011100000100011000011110000110100111101001001010001111000100011001001100011110100011010001111110010111000010110000111010010101000000001000110110001010100111000000100110010110100000101000001010010100000010000001101000001000100111100;
		
		// 32, 64
		//points = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010001001010001001000110101000111000001010000101001000011110001001100111101001111000011011100000110000011100010110000011001000111010001000000101000001100000010011100011001001001010001111100100011001101110000010000011111000111110010000100110001000100010000110000010100001001110010010100111111001011100000111100110101000110010011000100110100000000100010100000001101000011110000101100011011000000010001100000001001000101000001111000111101000110110010001100010011001111000011111000000011001100000001000100011100;
		
		// 64, 64
		//points = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001110000010101000111000010000000010010000110100010100000001101001101100000110000110011001001000010010000100111000000100000011100101101001000000010010000011110000101100011010100001000000100110001101000001110000001010000101000101101000011010010110000110101001110100000011100100111001000010010101100000000000011100011011000101010000101010001000000101111001101010011111000010100001011010001011000010100000100010011010000000111000100110001010100001001001110000011110000101001001100110000101100100101000000100001001100011111001111100000000000011011001111110011111100100111000110010001010000100101001101110001111100111100001011110011000000111100000000110000001000111111001111100000001000111111001110100010111100110100000011010000110100000110001110010011010100101011000010000010010000111100000001010001100100111011000110100011000100000110000101100000011100100110000010000001111000011001001010000001010000011000001100100000110100011000001111000010000100011100001100010010100100001111001010010011011100111110001010000000100100100010;
		
		// 256, 64
		points = 4096'b0001011000110011000111000010101000100101001000100001010000001011000111100011001000101100000010100001001100111101000000100000110100000001001010110010000100000011001110100010001100011111000100010001010100000001000110010000110000100010000111010001101000101110001111100010011100111110001001100001110000110111001110000011101100110111001011110000011000011110001111010000111100001001000001100011010100001011000101100000000000001011001000110010110000011111001100100000100000011010000111010001100100101101001100110010101100110001001011100011110000111110001011110010101000010111001001100011010100111111000100100010001100011011000011010001010100010111000001010011010100001011000011010011100000100011001000000011001000011000000001010000000100100101001110100011001000101010001111010001011100010010001101000001011100111101000010000001000000101100001000010010100000011010000111110001011100001000000010110011101000010111000011010010001100101101001010110010111000011100000010110001011100110011001101110000110000110111000101100001011000000011000010100000100000010110000000110001011100011011001001110010110100101100001001000001100000101100001010000001010000011001000101010000110000100011000101100010101100001001001100000011000100101010001110110000001100111111000000110011011100111011001110010001011100110000001111100011001000101011001101000000010000000001000110110000001100001010001110000011011000001001000000010001100000110000000101000010101100101100000100010001011000110111000001000001111000011010000110000010011000111110000011100001011100110111000011010010111000100100000010100010001100100110001000100011111100111111001010010000001100111010000110110011010100011000001100010010001100000000001010010000001100100111001011100000000000000111001000110000111000001000001111110011011000011110000100000011001100110110001110000010111000110101000010000010001000000010001011110000001000010111001001110000000000010110000001100010111000110001001110010010011100111111000100110011001100110010001111100001110100001011001011100000010000000001001111010001001000011111000010110001111000110111001100100010101000100000001000000001110000101100001101110000001000000110001000000001100000011001001101010010111100011110000011110010001000011100000101110001110000101110001011010000101100001110000100010011111000101111001010010000001100110001000000010011000000100100001011010001110100100100001000010000101000010100000100010011001100011011000000000011110100111010001110110010011000100100001011100011110000110111001101010001110000110011000101110010001000101000000100110000100100110100001101110010110000100001001111000010011000000111000010100011011100010001001001000000011100000000001010010000110000101000001111000000101000010011001011110000111100100010001110100000000000010010001001100010100100001101001111000001000000100010000111100000000000100101000111010000001000011010000111110010010000101001000001100011111100010110001100100010011000101100000100100001110000000000000111100000001000000111000000110010011100011100000110010001011000111010000100110000101100110011000111000010110000110010000101000010000100100011001010100001010000110100000010010011101100011001000000010011000000011000000000010001101100011011000001110010010100111111001001010000101100000100000101010001100000100101001000110011111100000101001110110010101100010001001100010010110100110010000100000000100100011011001010010010010100000010000111110010000100000010000101000000001000111100001101100011110100110011001111100010110100100001000100100010000100011000000000110001001100110110000100010001001000100000000011100010010000010000000111100010100000001001000101100001011100110101000000100011000000010100001101000001001100101001000101110011100100001001000110110011100000001100001010000000011100010111000101000001010000011111000101000010010100110010001011010001100000010011001111110010100100010111001100100010000100001001000011110001000100010100000111010010111100000001000010010011101000000100001001010011100000101010000100110001111100111100000111000000011100110101000101110000000000011101001001010000110100110100000111010011010100100011001111000001011000100101001110010000010000101110;
		
		// Wait for global reset to finish
		#100;
				
		// Generate a reset
		CPU_RESETN = 0;	#20;
		CPU_RESETN = 1;	#20;
		
		// Give a long time for machine to finish
		//#8000;
		//32000;
		#500000;
		
		// Wait for global reset to finish
		#100;

	end
		  
endmodule

