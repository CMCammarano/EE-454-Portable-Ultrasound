`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   20:12:24 10/05/2015
// Design Name:   quickhull.v
// 
////////////////////////////////////////////////////////////////////////////////

module m_quickhull_tb;

	// Inputs
	reg CLK100MHZ;
	reg CPU_RESETN;
	reg [4095:0] points;
	reg [7:0] SS;

	// Outputs
	wire [4095:0] convexPoints;
	wire [7:0] convexSetSize;
	wire [7:0] positiveCrossCount;
	wire [15:0] crossValue;
	wire [15:0] lnIndex;
	wire [7:0] ptCount;
	wire [31:0] currLine;
	wire [15:0] currPoint;
	wire [15:0] furthest;

	wire QINITIAL, QFIND_MAX, QFIND_MIN, QHULL_START, QCROSS, QHULL_RECURSE, QEND;
	// File
	integer file_results;

	// Parameters
	parameter CLK_PERIOD = 20;

	// Instantiate the Unit Under Test (UUT)
	m_port_ultra_quickhull_processor UUT(
		//Inputs
		.CLK100MHZ(CLK100MHZ),
		.CPU_RESETN(CPU_RESETN),
		.SS(SS),
		.points(points),
		//Outputs
		.convexPoints(convexPoints),
		.convexSetSizeOutput(convexSetSize),
		.positiveCrossCountOutput(positiveCrossCount),
		.crossValueOutput(crossValue),
		.lnIndexOutput(lnIndex),
		.ptCountOutput(ptCount),
		.currentLineOutput(currLine),
		.currentPointOutput(currPoint),
		.furthestOutput(furthest),
		.QINITIAL(QINITIAL),
		.QFIND_MAX(QFIND_MAX),
		.QFIND_MIN(QFIND_MIN),
		.QHULL_START(QHULL_START),
		.QCROSS(QCROSS),
		.QHULL_RECURSE(QHULL_RECURSE),
		.QEND(QEND)
	);


	initial begin : CLOCK_GENERATOR
		CLK100MHZ = 0;
		
		forever begin
			# (CLK_PERIOD / 2) CLK100MHZ = ~CLK100MHZ;
		end
	end	
		
	integer counter;
	
	initial begin : STIMULUS
		
		//file_results = $fopen("output_results.txt", "w");

		// Initialize Inputs
		// === Small input: 15 points ===
		/*
		SS = 15;
		
		points = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000011000000101000010000000001100000111000001110000100100000111000001000000001000000101000001010000000100000100000001100000010100000011000001000000001000000100000001010000010100000110000000110000010000001100000010010000101100000001;


		// Wait for global reset to finish
		#100;
				
		// Generate a reset
		CPU_RESETN = 0;	#20;
		CPU_RESETN = 1;	#20;
		
		// Give a long time for machine to finish
		#500000;

		//$fwrite(file_results, "Points:     ");
		$write("Points:     ");
		
		// Wait for global reset to finish
		#100;
		*/
		// === Medium input: 50 points ===
		//Input next test
		SS = 50;

		//Range: 0 - 31
		/*
		points = 4096'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001010000010000000011000000100000000000000111100010011000111110001101000010010000100010001110100011011000101100001011000010100000100100000011000011111000001110000010000010101000010010000101100001110000011000000010000011010000111100001011100000011000111000000110000001101000000110001011100001111000000010001111000000011000001000001111000010010000100000000111100010010000111110001101000000100000011000001111100000010000110100000011000011011000110110001101100011011000110000001001100000010000000110000001000011100000110100000111000001101000100110000011100001110000010110001000000010011000111010000011100011111000101000001001100010110000001000001111100000110000001000000111100011000000100000000000100001110000000010000100100010011000001010001111100010101000011110001110000000000000001100001010000001100;
		*/
		
		points = 0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100001011100100000110101110110001110000010101100111011011011100101011001111001011011010011001100110110011000000000101101001110000000110101101001010001001111010110100101100011000011110001010000010100010100110001101100111000010110110011100101010100001111110011111000011111010001000110010101111010000010010010100100101111001100100000011001111011011001010011011101101111010010110001011101001111010010010000101000000011001111010011111101100111000110000010111101010011001101000001101001000111010001010100000100110011010100110011100001000111001000010000100100000101001100000011000000010011001101010011111000100000001001110001010000100100011011100101110001010110010000110111001000011100011000100000110000000110011011010011000101100011010010000000000001010101010110010011101001110110001110100111010001111100001011000100011100001100000001010100011100100010010011010001011001010110001110100100010100110111001100000010010101011010000001100000011001011010000010100100000101100001000110010001101101000011010001110100110100111010011101110011110001011110010001100010110001100100001101100101100001001100000010110000101001101110011111000011011000110101010000000010011101011110011111100110101101100001000100110111111101000000011110010000110000101001001000110110000101100111011101000111001101000010000101010101111100100010000101000000101100001000011001100010010100000101001000010011011000100100000011110111110100100000001001100010101100000000010011010111000100001011010000000100100101100111010001000010110101011000000100000110000001101101011010110001010001000110001111100010010100000010011011000100010101101000001101100001100000010111011000010110001100000010010000100110000101001001001100010010100100110111010101110001010001100110010011110100111000011011000101000001011001011100001000100100100001111100010111100101011101010100011111000011111000000011001111010110100101011100001101100101001000011100011001110010001000110100000001110010111000001011001010110101101100000111000100110111010101010010001110000100110101000100000100100101011101101100011101100011101101110101;
		// Wait for global reset to finish
		#100;
				
		// Generate a reset
		CPU_RESETN = 0;	#20;
		CPU_RESETN = 1;	#20;
		
		// Give a long time for machine to finish
		#5000000;
		
		/*
		// === Max input: 256 points ===
		// Input next test
		SS = 255;

		//Range 0 - 31
		points = 4096b'0001110000010100000011010000101100010101000011010000011100010110000110110000001100001001000101000001111000011111000101000001011100011100000100010001000000010110000100000001011000011011000101010001000000010111000001000000010000000001000110010000111000000101000111000000000100010000000100010000101000001000000000110001110100001100000100100000110100001000000111010001111000000011000100110000101000001101000001110000001100010010000101000000101000010111000010100001101000000001000010110001001100000111000010000000110100000100000000100000111000011011000000110001110000011011000001100001110000000100000010100000110000001001000001110000001100011110000001010000000100011011000100000000110000010100000100010001000100011000000000000001101000010100000011100000011100000101000000100000000100010111000010010000111100001000000001000001001000010000000011110000100100001110000100110001110100001110000000000000100100010010000010010001100000011010000001010000110000000100000100100001001000000100000101000001111000001001000100100000001000011011000101110000010100000010000000000000010100001000000010100000000000010100000001010000110000000100000001100001110000000101000011000000010000010001000111000000110000011100000001100000001100001101000010100000001000000100000101110001100100000101000101000000011000001010000111100001001100001001000011100000110100011000000101010001101000000010000110110001101100011011000101010001000100010010000111010001101100010101000010100001111000001000000100010001110100000110000101100000100100011001000001110001100000011110000100010000111000000011000000010000111100011101000101100001011000011101000110010000010000001011000111010000010000000110000010010000111100001100000001110000101000000011000110110000100000000000000100100000001100011101000010110001000100010001000101100001010100011110000100000001111100000011000011100000000000001010000111000001101100001111000000000000110000000001000111110000001000010101000000010001000000001100000101100001100000010001000111100001001100000100000010010000001100000011000111100000110000001111000000110000111100010000000101100000011100010010000100000001110100000011000000000000110000010011000101010000110000011101000000010000010000000001000111000001011100000000000011000001000000010100000111110001110000011111000011100000101000010001000110010001110100001010000100100000110100000100000001010001101100011000000110100000110100000110000000010000111100001111000100100000101100001110000110110001011100010110000001100000111000001111000001010000100100001001000001100000110100011011000100110001001100001101000010110001110100001111000101000000101000011010000111010001111100010100000010010001010100000010000011110000010000011010000001000001110000010110000000110001010100010001000111110001001000010100000111110001001000010001000001100000011100001011000000110001101100010110000101100000110000001010000111010000101100000111000100000001110000010000000001110001110100010010000101110001101000011000000111110001000100010100000110010001111100000011000101100000100100000011000111010001011000011000000011100000010100001000000000010000000000001011000111100001011000000010000011100000011100010110000011000000011100010101000001010000001000001101000100100001010100011110000100000000110000001110000100010000001100011000000000100001100100011100000111000001101100001000000100100001101100001000000011000001100000010110000110100001110000000011000000110000001000000111000111110001001100011111000000100000101000010001000010110000110000011111000110110001000000000101000100110001011000000101000101110000010000011010000100000000111000011101000110010001010000001001000101000001010100011010000010110000001000010111000100000000111000011010000100000001101000001011000110000001111000001001000100000001001100010011000110100001011000010000000010100001011100001100000110110000110000010111000111000001001000001111000100110001111000011001000100110000110000010100000011000000110000000111000100100001111100001110000010110000001100010011000110100001111000001001000011010000010100010001000001010001011100000101000110100001000000011110000100100001111100001111000111100000100000000110000111000001001000000101;

		//Range 0 - 255
		//points =  4096'b0101110111110101111110100000100001100000111110100110001101001011011010000010110001110001100000011000011111001101011101100001010100010100000010111000111100011000101110101110011101000100101010110010100100010111100111000110011000010010000110010111111010000011000100000001110111101100001110001100001110000100010110111110100110011011011000000100010110001001001011100001111110100101101001101101000010010001011110001010100000100001010111011101110011000011001000001100011001111010111000110010000101111101110110110101000000011011001100100111110010101101100011111010010101001001010010110111011111100100100100001111110011111001100010000110100101100011101010001010001011000110010000010110101110001011011001001000100011100011000100110011000101111010010100010100101110100010011000111011011001011011011100000011010001100101110111101111111100101010101101001100011010111000100010101110101010111100111100000010011101101011101110000100011011011010110111000101100111100001111110101110000111010110111111011101010100100010011001010001111000110110010011110110010110000100001000010001110100110110111101000000000001011010110000111101100001111010000001100111111010101110111010110010110010110100110100010101000001010000011110001100101001010001011011100100110111001011010000100011001000001001000011101010010010100011010100001110100011100000000101101111000110000110000001000100100110000010010001100101000011001111011010110010111010100110111101000101000111101111001010010011101100110111010010111110001111011010000000010011111110100010100010010011010111010101101110000100000010110000111000110111000011111000001011001101100010110110100101010100111010110100000011010000100100110100101001100100010110101000010010110011111100011011110001001101001110001110000110011000001101001010011011011110000000100001001010100010001101100101111011110011001111001111001011110011110101001001011011011011111011110000100110011110101101010111010011101110011011101010111101110010111101110101110010011110001000000111010010100001110001001001010001010100110001110110001011010001110111110011000100111000110111001111100100111110000100000111000101110110111011110101100001000001011111000100001100000111010110000010010011011101100100111000001011011100011010111111001011010101101000011110000111100001001010010001111110011001111011111011001010111111111110111101101000100111110101011111111001000111110011000111110110000000101011010111101010101101101000111110100000000001101111100110101110011010001000111010010101110101101001010000011110111101000111000011000001110101100010100110001001000000100001010000010101110011011001110110011010100110001001000001001101010101111011110111011011011111111010110100011101011000000011010010001011100000000000100101000011101001010000000001110001101111100001000010100100001010111001010100010101100100101001111010010000000010011111000010101011101001111010011010110110100010101010100111011111001000101000010110100111000010000001010001011001011000100011111001010010000011100010001011001001100000110100001011000110100011001101000110110000001001101000101111111111011010101100101110111010111010001110001101001011110010111001000101100010000011101011110011001001100110011100001010000111100011001110001101101010011110100000100011100001101111101010101111110100101111100001110000101000001001111110010010101000000001010001001011111000011001110110010101001011000101101011100101110110111001110010110011000101000011001000110010001011110101000100110001110110011111001000111010111110001000010101111111010011111011111111010110001010000100011001101000011000111000110010010001100101011100001100100010011111100000111101110011101101100000000110110100001010111111010001011110011000101001011100001100001111001010010010001011000001000100101010011100010001101010001110001110000001010000100111011100111100100110101101001101111111010001110100100100001101101010111110000010011010010101010100010101011010111101010001100011001001111011010111110011110011110001110100110100001010111011000111011001101110100101111100001100100011001010111101111000001001000010110101010101110011000011101110001000110011100110001110101011110000001001100101100101010101011111110101011010;

		for (counter = 0; counter < convexSetSize; counter = counter + 1) begin
			//$fwrite(file_results, " %h", convexPoints[(16*counter)-1 +: (16*counter)]);
			//$write(file_results, " %h", convexPoints[(16*counter)-1 +: (16*counter)]);
		end


		// Wait for global reset to finish
		#100;
				
		// Generate a reset
		CPU_RESETN = 0;	#20;
		CPU_RESETN = 1;	#20;
		
		// Give a long time for machine to finish
		#10000;
		
		//$fwrite(file_results, "Points:     ");
		$write("Points:     ");
		*/
		// Wait for global reset to finish
		#100; 

	end
		  
endmodule

